library verilog;
use verilog.vl_types.all;
entity f1 is
end f1;
